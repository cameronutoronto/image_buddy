`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/24/2018 01:31:01 PM
// Design Name: 
// Module Name: slicer15
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module slicer15(
    input [14:0] din,
    output out00,
    output out01,
    output out02,
    output out03,
    output out04,
    output out05,
    output out06,
    output out07,
    output out08,
    output out09,
    output out10,
    output out11,
    output out12,
    output out13,
    output out14
    );
    
assign out00 = din[0];
assign out01 = din[1];
assign out02 = din[2];
assign out03 = din[3];
assign out04 = din[4];
assign out05 = din[5];
assign out06 = din[6];
assign out07 = din[7];
assign out08 = din[8];
assign out09 = din[9];
assign out10 = din[10];
assign out11 = din[11];
assign out12 = din[12];
assign out13 = din[13];
assign out14 = din[14];
endmodule
